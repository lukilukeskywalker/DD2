
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package Master_SPI_test_pack is

	constant Tclk_50_Mhz:	time:=20 ns;
