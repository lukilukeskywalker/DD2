--Autor LX0809 G4 Lukitas
